`timescale 1ns / 1ps

module hw2testbench(
    );

//wires
wire [16:0] finResult;

//regs
reg [15:0]x;
reg [15:0]y;
reg c16;
reg c;

top uut(
    .c(c),
    .x(x),
    .y(y),
    .c16(c16),
    .finResult(finResult)
);

initial begin
    c = 1'b0; //intialize the first carry value
    //Test Cases
    //15 + 1 = 16
    y = 16'b0000000000000010;
    x = 16'b0000000000001111;
    #2;
    y = 16'b000000000000001;
    x = 16'b000000000000001;
    #2;
    //3 + 3 = 6
    y = 16'b000000000000011;
    x = 16'b000000000000011;
    #2;
    //8 + 8 = 16
    y = 16'b000000000001000;
    x = 16'b000000000001000;
    #2;
    //15 + 15 = 30
    y = 16'b000000000001111;
    x = 16'b000000000001111;
    #2;
    //31 + 31 = 62
    y = 16'b000000000011111;
    x = 16'b000000000011111;
    #2;
    //12240 + 12901 = 135,301
    y = 16'd1224;
    x = 16'd12901;
    #2;
    //1224 + 32768 = 33,992
    y = 16'd12240;
    x = 16'd32768;
    #2;
    //66 + 400 = 466
    y = 16'd66;
    x = 16'd400;
    #2;
    //65535 + 400 == show over flow
    y = 16'b1111111111111111;
    x = 16'd600;
    #2;

end
endmodule